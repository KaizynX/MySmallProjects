`timescale 1ns / 1ps
module FullAdder();

endmodule // FullAdder