
module fdiv_s_p (
	source,
	probe);	

	output	[31:0]	source;
	input	[15:0]	probe;
endmodule
