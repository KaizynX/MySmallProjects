`timescale 1ns / 1ps
module FullAdder_Test();

FullAdder FA_Test();

endmodule // FullAdder_Test